
module mux4_32bit(sel, a0, a1, a2, a3, 
					which_a);
	input wire[1:0] sel;
	input wire[31:0] a0, a1, a2, a3;
	output wire[31:0] which_a;



endmodule // mux2_32bit
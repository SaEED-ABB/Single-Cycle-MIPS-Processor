
module sign_extend(a, 
					sign_extended_a);
	input wire[15:0] a;
	output wire[31:0] sign_extended_a;

	

endmodule // sign_extend

module instruction_memory(clk, rst, address, 
							instruction);
	input wire clk, rst;
	input wire[31:0] address;
	output wire[31:0] instruction;



endmodule // instruction_memory

module alu(ALUOperation, a, b, 
			zero, ALUResult);
	input wire[2:0] ALUOperation;
	input wire[31:0] a, b;
	output wire zero;
	output wire[31:0] ALUResult;
	
	
	
endmodule // alu

module shift_left2_32bit(a, 
						shifted_a);
	input wire[31:0] a;
	output wire[31:0] shifted_a;



endmodule // shift_left2_32bit 

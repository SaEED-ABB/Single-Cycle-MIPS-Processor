
module mux4_5bit(sel, a, b, c, d, 
					a_or_b_or_c_or_d);
	input wire[1:0] sel;
	input wire[4:0] a, b, c, d;
	output wire[4:0] a_or_b_or_c_or_d;

	

endmodule // mux2_32bit

module alu_control(clk, rst, instFunc, ALUOp, 
					ALUOperation);
	input wire clk, rst;
	input wire[5:0] instFunc;
	input wire[1:0] ALUOp;
	output wire[2:0] ALUOperation;



endmodule // alu_control

module shift_left16_16bit(a, 
						shifted_a);
	input wire[15:0] a;
	output wire[31:0] shifted_a;

	

endmodule // shift_left16_16bit
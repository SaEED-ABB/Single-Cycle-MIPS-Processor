
module pc_register(clk, rst, pc_in, 
					pc_out);
	input wire clk, rst;
	input wire[31:0] pc_in;
	output wire[31:0] pc_out;



endmodule // pc_register
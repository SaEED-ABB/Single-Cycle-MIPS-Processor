
module mux2_32bit(sel, a, b, 
					a_or_b);
	input wire sel;
	input wire[31:0] a, b;
	output wire[31:0] a_or_b;



endmodule // mux2_32bit